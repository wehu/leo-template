`include "leo_features.vh"

module dut(input int in, output int out);
  assign out = in;
endmodule
